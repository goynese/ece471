* # FILE NAME: /NFS/STAK/STUDENTS/G/GOYNESE/CADENCE/SIMULATION/LAB3CIRCUIT2/    
* HSPICES/SCHEMATIC/NETLIST/LAB3CIRCUIT2.C.RAW
* NETLIST OUTPUT FOR HSPICES.
* GENERATED ON JAN 31 16:21:29 2014
   
* GLOBAL NET DEFINITIONS
.GLOBAL VDD
* FILE NAME: ECE471_LAB3CIRCUIT2_SCHEMATIC.S.
* SUBCIRCUIT FOR CELL: LAB3CIRCUIT2.
* GENERATED FOR: HSPICES.
* GENERATED ON JAN 31 16:21:29 2014.
   
R0 NET6 NET06  400.0 M=1.0 
C3 NET06 0  500E-15 M=1.0 
C0 NET6 0  500E-15 M=1.0 
XI1 NET06 OUT INVERTER2_G1 
XI0 IN NET6 INVERTER2_G1 
   
   
   
   
* FILE NAME: ECE471_INVERTER2_SCHEMATIC.S.
* SUBCIRCUIT FOR CELL: INVERTER2.
* GENERATED FOR: HSPICES.
* GENERATED ON JAN 31 16:21:29 2014.
   
* TERMINAL MAPPING: IN = IN
*                   OUT = OUT
.SUBCKT INVERTER2_G1 IN OUT 
MN0 OUT IN 0 0  TSMC25DN  L=240E-9 W=480E-9 AD=288E-15 AS=288E-15 PD=2.16E-6 
+PS=2.16E-6 M=1 
MP0 OUT IN VDD VDD  TSMC25DP  L=240E-9 W=480E-9 AD=288E-15 AS=288E-15 
+PD=2.16E-6 PS=2.16E-6 M=1 
   
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS INVERTER2_G1 
   
.lib "/nfs/guille/u1/c/cdsmgr/cdsmgr/pdk/CDK1.4/local/models/hspice/public/publicModel/tsmc25dN" NMOS 
.lib "/nfs/guille/u1/c/cdsmgr/cdsmgr/pdk/CDK1.4/local/models/hspice/public/publicModel/tsmc25dP" PMOS 
   
* INCLUDE FILES
   
   
   
   
   
   
* END OF NETLIST
.TEMP    25.0000    
.OP
.save
.OPTION  INGOLD=2 ARTIST=2 PSF=2
+        PROBE=0
.END
