* # FILE NAME: /NFS/STAK/STUDENTS/G/GOYNESE/CADENCE/SIMULATION/NOR2/HSPICES/    
* SCHEMATIC/NETLIST/NOR2.C.RAW
* NETLIST OUTPUT FOR HSPICES.
* GENERATED ON JAN 31 12:22:50 2014
   
* GLOBAL NET DEFINITIONS
.GLOBAL VDD! 
* FILE NAME: ECE471_NOR2_SCHEMATIC.S.
* SUBCIRCUIT FOR CELL: NOR2.
* GENERATED FOR: HSPICES.
* GENERATED ON JAN 31 12:22:51 2014.
   
MN3 NET10 OUT 0 0  TSMC25DN  L=240E-9 W=480E-9 AD=288E-15 AS=288E-15 
+PD=2.16E-6 PS=2.16E-6 M=1 
MN2 NET10 OUT 0 0  TSMC25DN  L=240E-9 W=480E-9 AD=288E-15 AS=288E-15 
+PD=2.16E-6 PS=2.16E-6 M=1 
MN1 OUT NET39 0 0  TSMC25DN  L=240E-9 W=480E-9 AD=288E-15 AS=288E-15 
+PD=2.16E-6 PS=2.16E-6 M=1 
MN0 OUT NET41 0 0  TSMC25DN  L=240E-9 W=480E-9 AD=288E-15 AS=288E-15 
+PD=2.16E-6 PS=2.16E-6 M=1 
MP2 NET37 OUT VDD! VDD!  TSMC25DP  L=240E-9 W=960E-9 AD=576E-15 AS=576E-15 
+PD=3.12E-6 PS=3.12E-6 M=1 
MP1 OUT NET43 NET29 VDD!  TSMC25DP  L=240E-9 W=960E-9 AD=576E-15 AS=576E-15 
+PD=3.12E-6 PS=3.12E-6 M=1 
MP0 NET29 NET45 VDD! VDD!  TSMC25DP  L=240E-9 W=960E-9 AD=576E-15 AS=576E-15 
+PD=3.12E-6 PS=3.12E-6 M=1 
MP3 NET10 OUT NET37 VDD!  TSMC25DP  L=240E-9 W=960E-9 AD=576E-15 AS=576E-15 
+PD=3.12E-6 PS=3.12E-6 M=1 
V3 IN_B NET39 0
V2 IN_A NET41 0
V1 IN_B NET43 0
V0 IN_A NET45 0
   
   
   

* INCLUDE FILES
   
   
   

.END
