* # FILE NAME: /NFS/STAK/STUDENTS/G/GOYNESE/CADENCE/SIMULATION/LAB3CIRCUIT2/    
* HSPICES/EXTRACTED/NETLIST/LAB3CIRCUIT2.C.RAW
* NETLIST OUTPUT FOR HSPICES.
* GENERATED ON JAN 31 15:58:52 2014
   
* FILE NAME: ECE471_LAB3CIRCUIT2_EXTRACTED.S.
* SUBCIRCUIT FOR CELL: LAB3CIRCUIT2.
* GENERATED FOR: HSPICES.
* GENERATED ON JAN 31 15:58:52 2014.
   
C2 GND VDD  235.9049376E-15 M=1.0 
C3 GND 1  88.9994016E-15 M=1.0 
M4 OUT 1 VDD VDD  TSMC25DP  L=239.99999143598E-9 W=959.999965743918E-9 
+AD=576.000022418227E-15 AS=576.000022418227E-15 PD=2.15999989450211E-6 
+PS=2.15999989450211E-6 M=1 
M5 1 IN VDD VDD  TSMC25DP  L=239.99999143598E-9 W=959.999965743918E-9 
+AD=576.000022418227E-15 AS=576.000022418227E-15 PD=2.15999989450211E-6 
+PS=2.15999989450211E-6 M=1 
M6 OUT 1 GND GND  TSMC25DN  L=239.99999143598E-9 W=479.999982871959E-9 
+AD=288.000011209114E-15 AS=288.000011209114E-15 PD=1.67999996847357E-6 
+PS=1.67999996847357E-6 M=1 
M7 1 IN GND GND  TSMC25DN  L=239.99999143598E-9 W=479.999982871959E-9 
+AD=288.000011209114E-15 AS=288.000011209114E-15 PD=1.67999996847357E-6 
+PS=1.67999996847357E-6 M=1 
   
   
   
   
   
.lib "/nfs/guille/u1/c/cdsmgr/cdsmgr/pdk/CDK1.4/local/models/hspice/public/publicModel/tsmc25dN" NMOS 
.lib "/nfs/guille/u1/c/cdsmgr/cdsmgr/pdk/CDK1.4/local/models/hspice/public/publicModel/tsmc25dP" PMOS 
   
* INCLUDE FILES
   
   
   
   
   
   
* END OF NETLIST
.TEMP    25.0000    
.OP
.save
.OPTION  INGOLD=2 ARTIST=2 PSF=2
+        PROBE=0
.END
